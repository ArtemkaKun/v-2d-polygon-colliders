module pcoll2d
