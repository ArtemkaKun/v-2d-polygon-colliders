module pcoll2d

import artemkakun.trnsfrm2d

fn test_decompose_convex_polygon() {
	polygon := Polygon{
		points: [trnsfrm2d.Position{
			x: 0.0
			y: 0.0
		}, trnsfrm2d.Position{
			x: 0.0
			y: 1.0
		}, trnsfrm2d.Position{
			x: 1.0
			y: 1.0
		}, trnsfrm2d.Position{
			x: 1.0
			y: 0.0
		}]
	}
}
