module pcoll2d

fn decompose(polygon_points Polygon) []Polygon {
}
